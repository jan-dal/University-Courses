2b 5b 2d 5b 3c 3c 5b 2b 5b 2d 2d 2d 3e 5d 2d 5b 3c 3c 3c 5d 5d 5d 3e 3e 3e 2d 5d 3e 2d 2e 2d 2d 2d 2e 3e 2e 2e 3e 2e 3c 3c 3c 3c 2d 2e 3c 2b 2e 3e 3e 3e 3e 3e 2e 3e 2e 3c 3c 2e 3c 2d 2e 